'timescale 1ns/1ps

module echo_tx_ctrl (
    input wire  sys_clk    ,
    input wire  sys_rst    ,
    input wire [63:0]  echo_tx_data   ,
    input wire         echo_tx_en     ,
    output wire [63:0]  srio_tx_data    ,
    output wire         srio_tx_en    
);


endmoudle
